----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:25:44 10/24/2013 
-- Design Name: 
-- Module Name:    Hazarddetection - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Hazarddetection is
    Port ( IDEXCONTROL : in  STD_LOGIC_VECTOR(8 downto 0);
           IDEXregisterRT : in  STD_LOGIC_VECTOR(4 downto 0);
			  IFIDregisterRS : in  STD_LOGIC_VECTOR(4 downto 0);
			  IFIDregisterRT : in  STD_LOGIC_VECTOR(4 downto 0);
			  IFIDInstructionType: in  STD_LOGIC_VECTOR (5 downto 0);
           PCWrite : out  STD_LOGIC;
			  IFIDwrite: out STD_LOGIC;
			  IFIDreset: out STD_LOGIC;--remove this maybe?
			  processor_enable: in std_logic;
           Controlenable : out  STD_LOGIC

			  );
end Hazarddetection;



architecture Behavioral of Hazarddetection is


begin
	

process(processor_enable,IDEXCONTROL,IDEXregisterRT,IFIDregisterRS,IFIDregisterRT,IFIDInstructionType)
constant LW  : std_logic_vector(8 downto 0 ) := "000001110";
constant load  : std_logic_vector(5 downto 0 ) := "100011";
    constant BEQ  : std_logic_vector(5 downto 0 ) := "000100";
	 constant BNE  : std_logic_vector(5 downto 0 ) := "000101";
	 	 constant branchne  : std_logic_vector(8 downto 0 ) := "001-10000";
	 constant branche  : std_logic_vector(8 downto 0 ) := "101-00000";
begin


        if(processor_enable='1') then  
				
				if(IDEXCONTROL=LW and (IDEXregisterRT = IFIDregisterRS or IDEXregisterRT=IFIDregisterRT) AND NOT (IFIDInstructionType=LOAD)) then
				pcWrite<='0';
				ifidwrite<='0';
				Controlenable<='0';
				elsif (((IFIDInstructionType=BEQ) or (IFIDInstructionType=BNE)))then --and not( IDEXCONTROL=Branche or IDEXCONTROL=branchne)) then
				pcWrite<='0';
				ifidwrite<='1';
				Controlenable<='1';
				else
				pcWrite<='1';
				ifidwrite<='1';
				Controlenable<='1';
				end if;
				else
				PCWrite<='0';
				Controlenable<='0';
				ifidwrite<='1';
				
				end if;
end process;


end Behavioral;

