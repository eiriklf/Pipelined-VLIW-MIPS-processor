--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 


library IEEE;
use IEEE.STD_LOGIC_1164.all;

package Customtype is

  

type ProOP is (jump,memwrite,regwrite,memtoreg,alusrc,branch,regdest);


-- Declare constants


 

 
end Customtype;
